// file: InstMem.v
// author: @hazemwalidf

`timescale 1ns/1ns

module InstMem (
input [5:0] addr, 
output [31:0] data_out
    );
    reg [31:0] mem [0:63];
    assign data_out = mem[addr];
    
 initial begin
 
     mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
     //added to be skipped since PC starts with 4 after reset
     mem[1]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
     mem[2]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
     mem[3]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
     // mem[4]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
     mem[4]=32'b000000001001_00001_110_00100_0010011 ; //ori x4, x1, 9
     // mem[5]=32'b0_000000_00011_00100_000_0100_0_1100011; //beq x4, x3, 4
     // mem[5]=32'b0_000000_00010_00001_001_0100_0_1100011; //bne x1, x2, 4
     // mem[5]=32'b0_000000_00001_00010_100_0100_0_1100011; //blt x2, x1, 4
     // mem[5]=32'b0_000000_00010_00001_101_0100_0_1100011; //bge x1, x2, 4
     // mem[5]=32'b0_000000_00001_00010_110_0100_0_1100011; //bltu x2, x1, 4
     mem[5]=32'b0_000000_00010_00001_111_0100_0_1100011; //bgeu x1, x2, 4
     mem[6]=32'b0000000_00010_00001_100_00011_0110011 ; //add x3, x1, x2     
     // mem[7]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
     mem[7]=32'b000000001001_00011_000_00101_0010011 ; //addi x5, x3, 9
     mem[8]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
     mem[9]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
     // mem[10]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
     mem[10]=32'b000000111111_00110_111_00111_0010011 ; //andi x7, x6, 63
     mem[11]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
     mem[12]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
     mem[13]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
     mem[14]=32'b000000000101_00010_100_01010_0010011 ; //xori x10, x2, 5
     mem[15]=32'b0000000_00001_00010_001_01011_0010011 ; //slli x11, x2, 1
     mem[16]=32'b0000000_00001_01011_101_01100_0010011 ; //srli x12, x11, 1
     mem[17]=32'b0100000_00001_01011_101_01101_0010011 ; //srai x13, x11, 1
     mem[18]=32'b000000000010_00000_000_01110_0010011 ; //addi x14, x0, 2
     mem[19]=32'b0000000_01110_00010_001_01111_0110011 ; //sll x15, x2, x14 
     mem[20]=32'b0000000_01110_01111_101_10000_0110011 ;  //srl x16, x15, x14
     mem[21]=32'b000000001010_00010_010_10001_0010011 ; //slti x17, x2, 10
     mem[22]=32'b0000000_00001_00010_010_10010_0110011 ; //slt x18, x2, x1
     mem[23]=32'b0000001_01001_01001_000_10011_0110011 ; //mul x19, x9, x9
     mem[24]=32'b111111111110_00000_000_10100_0010011 ; //addi x20, x0, -2
     mem[25]=32'b0000001_10100_00001_001_10101_0110011 ; //mulh x21, x1, x20
     mem[26]=32'b0000001_00001_10100_010_10110_0110011 ; //mulhsu x22, x1, x20
     mem[27]=32'b0000001_01110_01001_110_10111_0110011 ; //rem x23, x9, x14
     
     
    // mem[23]=32'b0_0000001010_0_00000000_10011_1101111 ; //jal x19, 20
    // mem[24]=32'b000000001000_10000_000_10100_1100111 ; //jalr x20, 0(x19)
     
     
     /*
     mem[0]=32'h00400093;      //addi x1,x0,4 #x1=4                        
     mem[1]=32'h00800113  ;    //addi x2,x0,8 #x2=8                        
     mem[2]=32'h00300193  ;    //addi x3,x0,3 #x2=3                        
     mem[3]=32'h21100213  ;    //addi x4,x0,529 #x4=529                     
     mem[4]=32'h0010a023  ;    //sw x1,0(x1) # mem(4)=4                    
     mem[5]=32'h00412023  ;    //sw x4,0(x2) # mem(8)=528                  
     mem[6]=32'h00410223  ;    //sb x4,4(x2) # mem(12)=528                  
     mem[7]=32'h001102a3  ;    //sb x1,5(x2) # mem(13)=4                    
     mem[8]=32'h00411423  ;    //sh x4,8(x2) # mem(13)=528                  
     mem[9]=32'h00111523  ;    //sh x1,10(x2) # mem(13)=100                 
     mem[10]=32'h00012503 ;    //lw x10,0(x2) # x10= 528                   
     mem[11]=32'h00510583 ;    //lb x11,5(x2) # x11= 4 
     mem[12]=32'b0000000_00010_01100_001_01010_0100011 ; // lh x12, 10(x2)
     */
     
end



endmodule